�+�l�~���,r���O�@w?    ��?  �?                                          \
�b��b�W��9��O)q?    ��?  �?    �                                     ��ö���׵3��;뿱�>ԭ>   @��L?��L�    �                                     �[i����Sj�5;���=�[��=   @��L?��L�    �                                     �3��g?o�CښA���>   @��L?��L�                  8N�h����<��C,�       �/�擿�p|ÿ!���8?   @��L?��L�    �              �kk@ni���jB#��       *�H����<���?�H���>   @��L?��L�    @              A�+A�ٿ}H�u�˿       �j��c��f(�V���?׏�C�>   @��L?��L�    `	              A�+A�ٿ}H�u�˿       �>꧱a����ȁ���?�h��8>   @��L?��L�    �              A�+A�ٿ}H�u�˿       ��:��a���K�����?o����=   @��L?��L�    �              A�+A�ٿ}H�u�˿       鐲��a��������?.3�%7r=   @��L?��L�    �              A�+A�ٿ}H�u�˿       e�ٳ��?�{+�fN�?��y|[�?   @��L?��L�    x              E},��޿�r �I���       ����v��q��tr�ĿpW�Lΰ�>   @��L?��L�    (
              E},��޿�r �I���       H�3�_v��c6}�7�Ŀ��#��+>   @��L?��L�    �              E},��޿�r �I���       H�%�v�M���G�ܿN�1.��?   @��L?��L�    �              ����@ܿ45��Aܿ       \�!�3����Q^��ſG������>   @��L?��L�    �                                     5�� {�����E7
��m
�}]�>   @��L?��L�    (
                                     