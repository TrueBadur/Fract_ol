��ö���׵3��;뿱�>ԭ>   @��L?��L�    �                                     �[i����Sj�5;���=�[��=   @��L?��L�    �                                     �/�擿�p|ÿ!���8?   @��L?��L�    �              �kk@ni���jB#��       *�H����<���?�H���>   @��L?��L�    @              A�+A�ٿ}H�u�˿       �j��c��f(�V���?׏�C�>   @��L?��L�    `	              A�+A�ٿ}H�u�˿       �>꧱a����ȁ���?�h��8>   @��L?��L�    �              A�+A�ٿ}H�u�˿       ��:��a���K�����?o����=   @��L?��L�    �              A�+A�ٿ}H�u�˿       e�ٳ��?�{+�fN�?��y|[�?   @��L?��L�    x              E},��޿�r �I���       ����v��q��tr�ĿpW�Lΰ�>   @��L?��L�    (
              E},��޿�r �I���       H�3�_v��c6}�7�Ŀ��#��+>   @��L?��L�    �              E},��޿�r �I���       H�%�v�M���G�ܿN�1.��?   @��L?��L�    �              ����@ܿ45��Aܿ       \�!�3����Q^��ſG������>   @��L?��L�    �                                     5�� {�����E7
��m
�}]�>   @��L?��L�    (
                                     J8�����+\|O%7�?p�ds�>~�@�1M?��L�    d       ����    5��bS�@"��'���?       ��4����?��u_�XZ�5��I?~�@�1M?��L�                   �\����@a�䧂&��       ��V���"!�1��?���'�A?~�@�1M?��L�                   �>fOH��ߔ�Ț?       |8����?�h��->ſ��Gf���>      ��   @    @              ���WX��=h8�?       �2]B��ĸ�$x�ؿ -�:�=      ��   @    �                                     ��(�K��;d���V׿�e�5�>�ߔ�?�п���    �                                     �cY ��� �a�:�"�!�t)7>   @��L?��L�    �                                     |8����?�h��->ſ��Gf���>�"�?�U@��տ    @              ���WX��=h8�?       �Y��Vw���i��`���w�I��~i=~�@�1M?��L�    �                                     $���^��{����?>��>,�=   @��L?��L�    �              A�+A�ٿ}H�u�˿       ����%L˿���Q�?�T��	>�� @t�M?��L�    �              <�������˚�~85��       